/*
 *		テスト用プラットフォームのコンポーネント記述ファイル
 *
 *  $Id$
 */

/*
 *  カーネルオブジェクトの定義
 */
import(<kernel.cdl>);

/*
 *  ターゲット非依存のセルタイプの定義
 */
import("syssvc/tSerialPort.cdl");
import("syssvc/tSysLog.cdl");
import("syssvc/tSysLogAdapter.cdl");
import("syssvc/tBanner.cdl");
import("syssvc/tTestService.cdl");
import("syssvc/tTestServiceAdapter.cdl");

/*
 *  ターゲット依存部の取り込み
 */
import("target.cdl");

/*
 *  システムログ機能のアダプタの組上げ記述
 */
cell tSysLogAdapter SysLogAdapter {
	cSysLog = rKernelDomain::SysLog.eSysLog;
};

/*
 *  テストプログラム用サービスのアダプタの組上げ記述
 */
cell tTestServiceAdapter TestServiceAdapter {
	cTestService = rKernelDomain::TestService.eTestService;
};

/*
 *  これ以降のセルは，カーネルドメイン内に含める
 */
region rKernelDomain {

/*
 *  システムログ機能の組上げ記述
 */
cell tSysLog SysLog {
	logBufferSize = 32;					/* ログバッファのサイズ */
	initLogMask = 0;					/* ログバッファに記録すべき重要度 */
	initLowMask = C_EXP("LOG_UPTO(LOG_DEBUG)");
									   	/* 低レベル出力すべき重要度 */
	/* 低レベル出力との結合 */
	cPutLog = PutLogTarget.ePutLog;
};

/*
 *  カーネル起動メッセージ出力の組上げ記述
 */
cell tBanner Banner {
	/* 属性の設定 */
	targetName      = BannerTargetName;
	copyrightNotice = BannerCopyrightNotice;
};

/*
 *  テストサービスの組上げ記述
 */
cell tTestService TestService {
	cSysLog = SysLog.eSysLog;
};
};
